interface class Observable;
    pure virtual function dispose subscribe(observer obs);
endclass : Observable
