interface class Observer;
    pure virtual function invoke();
endclass : Observer
