interface class Data;
    pure virtual function bit[7:0] getData();
endclass
