interface class Generator;
  pure virtual function Transaction getTransaction();
endclass
